module y86_computer_main();

endmodule
